module OR_struct(res, A, B);
input A, B;
output res;
or(res, A, B);
endmodule 