module AND_struct(res, A, B);
input A, B;
output res;
and(res, A, B);
endmodule 
