module AND_DF(res, A, B);
input A, B;
output res;
assign res = A & B;
endmodule 